/*
 * File: sim_top.sv
 * Project: new
 * Created Date: 29/04/2022
 * Author: Shun Suzuki
 * -----
 * Last Modified: 30/04/2022
 * Modified By: Shun Suzuki (suzuki@hapis.k.u-tokyo.ac.jp)
 * -----
 * Copyright (c) 2022 Hapis Lab. All rights reserved.
 * 
 */

`timescale 1ns / 1ps
module sim_top();

endmodule
